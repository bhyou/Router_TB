interface line_serial_inf #( nodes=300 )( input clk, input reset);

  :wq




endinterface
