class flit_t #(int TYPE_WIDTH=2,int DATA_WIDTH=32);
        bit [TYPE_WIDTH-1:0] ftype;
        bit [DATA_WIDTH-1:0] content;
endclass
