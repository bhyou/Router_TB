package noc_router_pkg;
        
  import serial_pkg::*;
  import router_pkg::*;
  
  `include "router_env.svh"
  
endpackage
