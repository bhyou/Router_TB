interface line_para_inf(

);

  



endinterface
